library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;


entity DeBounce is
    port(   CLK : in std_logic;
            Reset : in std_logic;
            BUTTON : in std_logic;
            RESULT : out std_logic
        );
end DeBounce;

architecture behav of DeBounce is

--the below constants decide the working parameters.
--the higher this is, the more longer time the user has to press the button.
constant COUNT_MAX : integer := 100000; 
--set it '1' if the button creates a high pulse when its pressed, otherwise '0'.
constant BTN_ACTIVE : std_logic := '1';

signal count : integer := 0;
type state_type is (idle,wait_time); --state machine
signal state : state_type := idle;

begin
  
process(Reset,CLK)
begin
    if(Reset = '1') then
        state <= idle;
        RESULT <= '0';
   elsif(rising_edge(CLK)) then
        case (state) is
            when idle =>
                if(BUTTON = BTN_ACTIVE) then  
                    state <= wait_time;
                else
                    state <= idle; --wait until button is pressed.
                end if;
                RESULT <= '0';
            when wait_time =>
                if(count = COUNT_MAX) then
                    count <= 0;
                    if(BUTTON = BTN_ACTIVE) then
                        RESULT <= '1';
                    end if;
                    state <= idle;  
                else
                    count <= count + 1;
                end if; 
        end case;       
    end if;        
end process;                  
                                                                                
end architecture behav;